`timescale 1ns / 1ps

`ifndef _globals_vh_
`define _globals_vh_

`define CLK_FREQ 50_000_000

`endif
